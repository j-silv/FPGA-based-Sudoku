--parallel in, parallel out 8-stage 8-bit shift register
--data is parallel shifted from the bottom to the top
--the first row LED segment data is shifted through to the last stage shift register
--the last stage shift register will be thus connected to the first row of the LED matrix
library ieee;
use ieee.std_logic_1164.all;

--package for 8-stage 8-bit shift register array type
package shift_register_array is
	type shift_register is array (8 downto 0) of std_logic_vector(7 downto 0);
end package shift_register_array;

library ieee;
use ieee.std_logic_1164.all;
library work;
use work.shift_register_array.all;

entity shift_stage is
	port(
		--if shift_en = '1', parallel shifting is enabled
		--if shift_out = '1', output rows are updated
		clk, shift_out, shift_en, rst :  in std_logic;
	
		--this is where the data will come in
		data_in : in std_logic_vector(7 downto 0);
		
		--this array corresponds to each row connected to the LED matrix
		row : out shift_register := (others => (others => '0'))
	);
end entity shift_stage;

architecture logic of shift_stage is
	--internally shifting data
	signal temp_row : shift_register := (others => (others => '0'));
begin
	process(rst,clk)
	begin 
		if rst ='1' then
			temp_row <= (others => (others => '0'));
		else 
			if rising_edge(clk) then
				--is shifting through the stages enabled?
				if shift_en = '1' then
					--parallel shift in the first row information
					temp_row(8) <= data_in;
					
					--iterate and shift data through each stage once
					for i in 0 to 7 loop
						temp_row(7-i) <= temp_row(8-i);	
					end loop;
				end if;
			end if;
		end if;
	end process;
	
	process(shift_out)
	begin
		if rising_edge(shift_out) then
			--update LED segment data for LED matrix
			row <= temp_row;
		end if;
	end process;
end architecture logic;